`define TEST_NAME_STRING "or1k"
`define MOR1KX_CPU_PIPELINE cappuccino
