////////////////////////////////////////////////////////////////////////////////
//                                            __ _      _     _               //
//                                           / _(_)    | |   | |              //
//                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              //
//               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              //
//              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              //
//               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              //
//                  | |                                                       //
//                  |_|                                                       //
//                                                                            //
//                                                                            //
//              MPSoC-OR1K CPU                                                //
//              Processing Unit                                               //
//              Wishbone Bus Interface                                        //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

/* Copyright (c) 2015-2016 by the author(s)
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 *
 * =============================================================================
 * Author(s):
 *   Paco Reina Campo <pacoreinacampo@queenfield.tech>
 */

module or1k_cache_lru #(
  parameter NUMWAYS = 2,

  // Triangular number
  parameter WIDTH = NUMWAYS*(NUMWAYS-1) >> 1
)
  (
    input      [WIDTH-1:0] current,
    output reg [WIDTH-1:0] update,

    input      [NUMWAYS-1:0] access,
    output reg [NUMWAYS-1:0] lru_pre,
    output reg [NUMWAYS-1:0] lru_post
  );

  reg [NUMWAYS-1:0] expand [0:NUMWAYS-1];

  integer i, j;
  integer offset;

  // <    0      1      2      3
  // 0    1    (0<1)  (0<2)  (0<3)
  // 1  (1<0)    1    (1<2)  (1<3)
  // 2  (2<0)  (2<1)    1    (2<3)
  // 3  (3<0)  (3<1)  (3<2)    1
  //
  // As two entries can never be equally old (needs to be avoided on
  // the outside) this is equivalent to:
  //
  // <    0      1      2      3
  // 0    1    (0<1)  (0<2)  (0<3)
  // 1 !(0<1)    1    (1<2)  (1<3)
  // 2 !(0<2) !(1<2)    1    (2<3)
  // 3 !(0<3) !(1<3) !(2<3)    1
  //
  // The lower half below the diagonal is the inverted mirror of the
  // upper half. The number of entries in each half is of course
  // equal to the width of our LRU vector and the upper half is
  // filled with the values from the vector.
  //
  // The algorithm works as follows:
  //
  //  1. Fill the matrix (expand) with the values. The entry (i,i) is
  //     statically one.
  //
  //  2. The LRU_pre vector is the vector of the ANDs of the each row.
  //
  //  3. Update the values with the access vector (if any) in the
  //     following way: If access[i] is set, the values in row i are
  //     set to 0. Similarly, the values in column i are set to 1.
  //
  //  4. The update vector of the lru history is then generated by
  //     copying the upper half of the matrix back.
  //
  //  5. The LRU_post vector is the vector of the ANDs of each row.
  //
  // In the following an example will be used to demonstrate the algorithm:
  //
  //  NUMWAYS = 4
  //  current = 6'b110100;
  //  access  = 4'b0010;
  //
  // This current history is:
  //
  //  0<1 0<2 0<3 1<2 1<3 2<3
  //   0   0   1   0   1   1
  //
  // and way 2 is accessed.
  //
  // The history of accesses is 3>0>1>2 and the expected result is an
  // update to 2>3>0>1 with LRU_pre=2 and LRU_post=1

  always @(*) begin : comb
    // The offset is used to transfer the flat history vector into
    // the upper half of the
    offset = 0;

    // 1. Fill the matrix (expand) with the values. The entry (i,i) is
    //    statically one.
    for (i = 0; i < NUMWAYS; i = i + 1) begin
      expand[i][i] = 1'b1;
      for (j = i + 1; j < NUMWAYS; j = j + 1) begin
        expand[i][j] = current[offset+j-i-1];
      end
      for (j = 0; j < i; j = j + 1) begin
        expand[i][j] = !expand[j][i];
      end
      offset = offset + NUMWAYS - i - 1;
    end

    // For the example expand is now:
    // <    0      1      2      3        0 1 2 3
    // 0    1    (0<1)  (0<2)  (0<3)    0 1 0 0 1
    // 1  (1<0)    1    (1<2)  (1<3) => 1 1 1 0 1
    // 2  (2<0)  (2<1)    1    (2<3)    2 1 1 1 1
    // 3  (3<0)  (3<1)  (3<2)    1      3 0 0 0 1

    //  2. The LRU_pre vector is the vector of the ANDs of the each
    //     row.
    for (i = 0; i < NUMWAYS; i = i + 1) begin
      lru_pre[i] = &expand[i];
    end

    // We derive why this is the case for the example here:
    // lru_pre[2] is high when the following condition holds:
    //
    //  (2<0) & (2<1) & (2<3).
    //
    // Applying the negation transform we get:
    //
    //  !(0<2) & !(1<2) & (2<3)
    //
    // and this is exactly row [2], so that here
    //
    // lru_pre[2] = &expand[2] = 1'b1;
    //
    // At this point you can also see why we initialize the diagonal
    // with 1.

    //  3. Update the values with the access vector (if any) in the
    //     following way: If access[i] is set, the values in row i
    //     are set to 0. Similarly, the values in column i are set
    //     to 1.
    for (i = 0; i < NUMWAYS; i = i + 1) begin
      if (access[i]) begin
        for (j = 0; j < NUMWAYS; j = j + 1) begin
          if (i != j) begin
            expand[i][j] = 1'b0;
          end
        end
        for (j = 0; j < NUMWAYS; j = j + 1) begin
          if (i != j) begin
            expand[j][i] = 1'b1;
          end
        end
      end
    end

    // Again this becomes obvious when you see what we do here.
    // Accessing way 2 leads means now
    //
    // (0<2) = (1<2) = (3<2) = 1, and
    // (2<0) = (2<1) = (2<3) = 0
    //
    // The matrix changes accordingly
    //
    //   0 1 2 3      0 1 2 3
    // 0 1 0 0 1    0 1 0 1 1
    // 1 1 1 0 1 => 1 1 1 1 1
    // 2 1 1 1 1    2 0 0 1 0
    // 3 0 0 0 1    3 0 0 1 1

    // 4. The update vector of the lru history is then generated by
    //    copying the upper half of the matrix back.
    offset = 0;
    for (i = 0; i < NUMWAYS; i = i + 1) begin
      for (j = i + 1; j < NUMWAYS; j = j + 1) begin
        update[offset+j-i-1] = expand[i][j];
      end
      offset = offset + NUMWAYS - i - 1;
    end

    // This is the opposite operation of step 1 and is clear now.
    // Update becomes:
    //
    //  update = 6'b011110
    //
    // This is translated to
    //
    //  0<1 0<2 0<3 1<2 1<3 2<3
    //   0   1   1   1   1   0
    //
    // which is: 2>3>0>1, which is what we expected.

    // 5. The LRU_post vector is the vector of the ANDs of each row.
    for (i = 0; i < NUMWAYS; i = i + 1) begin
      lru_post[i] = &expand[i];
    end

    // This final step is equal to step 2 and also clear now.
    //
    // lru_post[1] = &expand[1] = 1'b1;
    //
    // lru_post = 4'b0010 is what we expected.
  end
endmodule
